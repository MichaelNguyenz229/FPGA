library verilog;
use verilog.vl_types.all;
entity my_tb is
end my_tb;
