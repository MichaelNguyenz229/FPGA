module first_practice
(
    input [31:0] a,
    input [31:0] b,
  
    output [31:0] add_out
);

assign add_out = a + b;

endmodule

